LIBRARY IEEE;
USE ieee.std_logic_1164.all;
-------------------------------
ENTITY serial_converter IS
	GENERIC ( MAX_WIDTH		:	INTEGER	:= 280);
	PORT	  ( clk				:	IN STD_LOGIC;
				 rst				:	IN	STD_LOGIC;
				 ena_guardar	:	IN STD_LOGIC;
				 ena_desplazar	:	IN STD_LOGIC;
				 transmitir		:	IN	STD_LOGIC_VECTOR (31 DOWNTO 0);
				 dout 			:	OUT STD_LOGIC:='1');
END ENTITY;
--------------------------------
ARCHITECTURE rtl OF serial_converter IS
	SIGNAL buffer_s: STD_LOGIC_VECTOR(MAX_WIDTH-1 DOWNTO 0);
	SIGNAL d			: STD_LOGIC_VECTOR(MAX_WIDTH-1 DOWNTO 0);
BEGIN
	
	d(9) <= '1'; -- bit parada
	d(8) <= '0';
	d(7) <= '1';
	d(6) <= '0';
	d(5) <= '1'; ------ t
	d(4) <= '0';
	d(3) <= '1';
	d(2) <= '0';
	d(1) <= '0'; 
	d(0) <= '0'; -- bit inicio
	d(19) <= '1'; -- bit parada
	d(18) <= '0';
	d(17) <= '1';
	d(16) <= '0';
	d(15) <= '0'; ------ i
	d(14) <= '1';
	d(13) <= '0';
	d(12) <= '0';
	d(11) <= '1'; 
	d(10) <= '0'; -- bit inicio
	d(29) <= '1'; -- bit parada
	d(28) <= '0';
	d(27) <= '1';
	d(26) <= '0';
	d(25) <= '0'; ------ e
	d(24) <= '0';
	d(23) <= '1';
	d(22) <= '0';
	d(21) <= '1'; 
	d(20) <= '0'; -- bit inicio
	d(39) <= '1'; -- bit parada
	d(38) <= '0';
	d(37) <= '1';
	d(36) <= '0';
	d(35) <= '0'; ------ m
	d(34) <= '1';
	d(33) <= '1';
	d(32) <= '0';
	d(31) <= '1'; 
	d(30) <= '0'; -- bit inicio
	d(49) <= '1'; -- bit parada
	d(48) <= '0';
	d(47) <= '1';
	d(46) <= '0';
	d(45) <= '1'; ------ p
	d(44) <= '0';
	d(43) <= '0';
	d(42) <= '0';
	d(41) <= '0'; 
	d(40) <= '0'; -- bit inicio
	d(59) <= '1'; -- bit parada
	d(58) <= '0';
	d(57) <= '1';
	d(56) <= '0';
	d(55) <= '0'; ------ o
	d(54) <= '1';
	d(53) <= '1';
	d(52) <= '1';
	d(51) <= '1'; 
	d(50) <= '0'; -- bit inicio
	d(69) <= '1'; -- bit parada
	d(68) <= '0';
	d(67) <= '0';
	d(66) <= '1';
	d(65) <= '0';
	d(64) <= '0'; ----- espacio
	d(63) <= '0';
	d(62) <= '0';
	d(61) <= '0'; 
	d(60) <= '0'; -- bit inicio
	d(79) <= '1'; -- bit parada
	d(78) <= '0';
	d(77) <= '1';
	d(76) <= '0';
	d(75) <= '0'; ------ d
	d(74) <= '0';
	d(73) <= '1';
	d(72) <= '0';
	d(71) <= '0'; 
	d(70) <= '0'; -- bit inicio
	d(89) <= '1'; -- bit parada
	d(88) <= '0';
	d(87) <= '1';
	d(86) <= '0';
	d(85) <= '0'; ------ e
	d(84) <= '0';
	d(83) <= '1';
	d(82) <= '0';
	d(81) <= '1'; 
	d(80) <= '0'; -- bit inicio
	d(99) <= '1'; -- bit parada
	d(98) <= '0';
	d(97) <= '0';
	d(96) <= '1';
	d(95) <= '0';
	d(94) <= '0'; ----- espacio
	d(93) <= '0';
	d(92) <= '0';
	d(91) <= '0'; 
	d(90) <= '0'; -- bit inicio
	d(109) <= '1'; -- bit parada
	d(108) <= '0';
	d(107) <= '1';
	d(106) <= '0';
	d(105) <= '0'; ------ e
	d(104) <= '0';
	d(103) <= '1';
	d(102) <= '0';
	d(101) <= '1'; 
	d(100) <= '0'; -- bit inicio
	d(119) <= '1'; -- bit parada
	d(118) <= '0';
	d(117) <= '1';
	d(116) <= '0';
	d(115) <= '0'; ------ j
	d(114) <= '1';
	d(113) <= '0';
	d(112) <= '1';
	d(111) <= '0'; 
	d(110) <= '0'; -- bit inicio
	d(129) <= '1'; -- bit parada
	d(128) <= '0';
	d(127) <= '1';
	d(126) <= '0';
	d(125) <= '0'; ------ e
	d(124) <= '0';
	d(123) <= '1';
	d(122) <= '0';
	d(121) <= '1'; 
	d(120) <= '0'; -- bit inicio
	d(139) <= '1'; -- bit parada
	d(138) <= '0';
	d(137) <= '1';
	d(136) <= '0';
	d(135) <= '0'; ------ c
	d(134) <= '0';
	d(133) <= '0';
	d(132) <= '1';
	d(131) <= '1'; 
	d(130) <= '0'; -- bit inicio
	d(149) <= '1'; -- bit parada
	d(148) <= '0';
	d(147) <= '1';
	d(146) <= '0';
	d(145) <= '1'; ------ u
	d(144) <= '0';
	d(143) <= '1';
	d(142) <= '0';
	d(141) <= '1'; 
	d(140) <= '0'; -- bit inicio
	d(159) <= '1'; -- bit parada
	d(158) <= '0';
	d(157) <= '1';
	d(156) <= '0';
	d(155) <= '0'; ------ c
	d(154) <= '0';
	d(153) <= '0';
	d(152) <= '1';
	d(151) <= '1'; 
	d(150) <= '0'; -- bit inicio
	d(169) <= '1'; -- bit parada
	d(168) <= '0';
	d(167) <= '1';
	d(166) <= '0';
	d(165) <= '0'; ------ i
	d(164) <= '1';
	d(163) <= '0';
	d(162) <= '0';
	d(161) <= '1'; 
	d(160) <= '0'; -- bit inicio
	d(179) <= '1'; -- bit parada
	d(178) <= '0';
	d(177) <= '1';
	d(176) <= '0';
	d(175) <= '0'; ------ o
	d(174) <= '1';
	d(173) <= '1';
	d(172) <= '1';
	d(171) <= '1'; 
	d(170) <= '0'; -- bit inicio
	d(189) <= '1'; -- bit parada
	d(188) <= '0';
	d(187) <= '1';
	d(186) <= '0';
	d(185) <= '0'; ------ n
	d(184) <= '1';
	d(183) <= '1';
	d(182) <= '1';
	d(181) <= '0'; 
	d(180) <= '0'; -- bit inicio
	d(199) <= '1'; -- bit parada
	d(198) <= '0';
	d(197) <= '0';
	d(196) <= '1';
	d(195) <= '1';	------ dos puntos
	d(194) <= '1';
	d(193) <= '0';
	d(192) <= '1';
	d(191) <= '0'; 
	d(190) <= '0'; -- bit inicio
	d(209) <= '1'; -- bit parada
	d(208) <= '0';
	d(207) <= '0';
	d(206) <= '1';
	d(205) <= '0';
	d(204) <= '0'; ----- espacio
	d(203) <= '0';
	d(202) <= '0';
	d(201) <= '0'; 
	d(200) <= '0'; -- bit inicio
	d(219) <= '1'; -- bit parada
	d(218) <= transmitir(31);
	d(217) <= transmitir(30);
	d(216) <= transmitir(29);
	d(215) <= transmitir(28);
	d(214) <= transmitir(27);
	d(213) <= transmitir(26);
	d(212) <= transmitir(25);
	d(211) <= transmitir(24);
	d(210) <= '0';
	d(229) <= '1';
	d(228) <= transmitir(23);
	d(227) <= transmitir(22);
	d(226) <= transmitir(21);
	d(225) <= transmitir(20);
	d(224) <= transmitir(19);
	d(223) <= transmitir(18);
	d(222) <= transmitir(17);
	d(221) <= transmitir(16);
	d(220) <= '0';
	d(239) <= '1';
	d(238) <= '0';
	d(237) <= '0';
	d(236) <= '1';
	d(235) <= '0';
	d(234) <= '1';
	d(233) <= '1';
	d(232) <= '1';
	d(231) <= '0';
	d(230) <= '0';
	d(249) <= '1';
	d(248) <= transmitir(15);
	d(247) <= transmitir(14);
	d(246) <= transmitir(13);
	d(245) <= transmitir(12);
	d(244) <= transmitir(11);
	d(243) <= transmitir(10);
	d(242) <= transmitir(9);
	d(241) <= transmitir(8);
	d(240) <= '0';
	d(259) <= '1';
	d(258) <= transmitir(7);
	d(257) <= transmitir(6);
	d(256) <= transmitir(5);
	d(255) <= transmitir(4);
	d(254) <= transmitir(3);
	d(253) <= transmitir(2);
	d(252) <= transmitir(1);
	d(251) <= transmitir(0);
	d(250) <= '0';
	d(269) <= '1';
	d(268) <= '0';
	d(267) <= '0';
	d(266) <= '1';
	d(265) <= '0';
	d(264) <= '0';
	d(263) <= '0';
	d(262) <= '0';
	d(261) <= '0';
	d(260) <= '0';
	d(279) <= '1';
	d(278) <= '0';
	d(277) <= '1';
	d(276) <= '1';
	d(275) <= '1';
	d(274) <= '0';
	d(273) <= '0';
	d(272) <= '1';
	d(271) <= '1';
	d(270) <= '0';
	PROCESS (clk, rst)
	BEGIN
		IF (rst='1') THEN
			buffer_s <= (OTHERS => '1');
		ELSIF (rising_edge(clk)) THEN
			IF (ena_guardar='1' AND ena_desplazar='0') THEN
				buffer_s <= d;
			ELSIF (ena_guardar='0' AND ena_desplazar='1') THEN
				buffer_s <= '1' & buffer_s(MAX_WIDTH-1 DOWNTO 1);
			ELSE
			buffer_s<= buffer_s;
			END IF;
		END IF;
	END PROCESS;
	
	dout <= buffer_s(0);
END ARCHITECTURE;