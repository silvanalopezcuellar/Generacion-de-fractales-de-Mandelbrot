LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--USE IEEE.STD_LOGIC_ARITH.ALL;
-------------------------
ENTITY register_cy0 IS
	GENERIC( DATA_WIDTH		:	INTEGER:= 32;
				ADDR_WIDTH		:	INTEGER);
	PORT(		clk				:	IN		STD_LOGIC;
				r_addr			:	IN		INTEGER;
				r_data			:	OUT	SIGNED(DATA_WIDTH-1 DOWNTO 0)				
			);
END ENTITY;
--------------------------
ARCHITECTURE rtl OF register_cy0 IS
	TYPE mem_2d_type IS ARRAY (0 TO ADDR_WIDTH) OF SIGNED((DATA_WIDTH)-1 DOWNTO 0);
	SIGNAL array_reg: mem_2d_type;
BEGIN
	--WRITE PROCESS
	array_reg(0)<= "11111100000000000000000000000000";
	
	array_reg(1)<= "00000000000000000000000000000000";
	array_reg(2)<= "00000000000000000000000000000000";
	array_reg(3)<= "11111100000000000000000000000000";
	array_reg(4)<= "11111100000000000000000000000000";
	
	array_reg(5)<= "00000010000000000000000000000000";
	array_reg(6)<= "00000010000000000000000000000000";
	array_reg(7)<= "00000000000000000000000000000000";
	array_reg(8)<= "00000000000000000000000000000000";
	
	array_reg(9)<= "00000010000000000000000000000000";
	array_reg(10)<= "00000010000000000000000000000000";
	array_reg(11)<= "00000000000000000000000000000000";
	array_reg(12)<= "00000000000000000000000000000000";
	
	array_reg(13)<= "11111110000000000000000000000000";
	array_reg(14)<= "11111110000000000000000000000000";
	array_reg(15)<= "11111100000000000000000000000000";
	array_reg(16)<= "11111100000000000000000000000000";
	
	array_reg(17)<= "11111110000000000000000000000000";
	array_reg(18)<= "11111110000000000000000000000000";
	array_reg(19)<= "11111100000000000000000000000000";
	array_reg(20)<= "11111100000000000000000000000000";
	
	--READ
	r_data <= array_reg(r_addr);
END ARCHITECTURE;